LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_unsigned.all;
USE ieee.std_logic_misc.all;
USE ieee.numeric_std.all;

-- ******************************************************************************
-- * License Agreement                                                          *
-- *                                                                            *
-- * Copyright (c) 1991-2013 Altera Corporation, San Jose, California, USA.     *
-- * All rights reserved.                                                       *
-- *                                                                            *
-- * Any megafunction design, and related net list (encrypted or decrypted),    *
-- *  support information, device programming or simulation file, and any other *
-- *  associated documentation or information provided by Altera or a partner   *
-- *  under Altera's Megafunction Partnership Program may be used only to       *
-- *  program PLD devices (but not masked PLD devices) from Altera.  Any other  *
-- *  use of such megafunction design, net list, support information, device    *
-- *  programming or simulation file, or any other related documentation or     *
-- *  information is prohibited for any other purpose, including, but not       *
-- *  limited to modification, reverse engineering, de-compiling, or use with   *
-- *  any other silicon devices, unless such use is explicitly licensed under   *
-- *  a separate agreement with Altera or a megafunction partner.  Title to     *
-- *  the intellectual property, including patents, copyrights, trademarks,     *
-- *  trade secrets, or maskworks, embodied in any such megafunction design,    *
-- *  net list, support information, device programming or simulation file, or  *
-- *  any other related documentation or information provided by Altera or a    *
-- *  megafunction partner, remains with Altera, the megafunction partner, or   *
-- *  their respective licensors.  No other licenses, including any licenses    *
-- *  needed under any third party's intellectual property, are provided herein.*
-- *  Copying or modifying any file, or portion thereof, to which this notice   *
-- *  is attached violates this copyright.                                      *
-- *                                                                            *
-- * THIS FILE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR    *
-- * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,   *
-- * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL    *
-- * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER *
-- * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING    *
-- * FROM, OUT OF OR IN CONNECTION WITH THIS FILE OR THE USE OR OTHER DEALINGS  *
-- * IN THIS FILE.                                                              *
-- *                                                                            *
-- * This agreement shall be governed in all respects by the laws of the State  *
-- *  of California and by the laws of the United States of America.            *
-- *                                                                            *
-- ******************************************************************************

-- ******************************************************************************
-- *                                                                            *
-- * This module connects the Avalon Switch Frabic to an External Bus           *
-- *                                                                            *
-- ******************************************************************************

ENTITY nios_system_to_external_bus_bridge_0 IS


-- *****************************************************************************
-- *                             Generic Declarations                          *
-- *****************************************************************************
	
GENERIC (
	
	AW		:INTEGER									:= 14;	-- Address bits
	EAB	:INTEGER									:= 1;		-- Extra address bits needed for the output address
	OW		:INTEGER									:= 15;	-- Address bits of the output port
	
	DW		:INTEGER									:= 15;	-- Data bits
	BW		:INTEGER									:= 1	--  Byte enable bits
	
);
-- *****************************************************************************
-- *                             Port Declarations                             *
-- *****************************************************************************
PORT (
	-- Inputs
	clk						:IN		STD_LOGIC;
	reset						:IN		STD_LOGIC;

	avalon_address			:IN		STD_LOGIC_VECTOR(AW DOWNTO  0);	
	avalon_byteenable		:IN		STD_LOGIC_VECTOR(BW DOWNTO  0);	
	avalon_chipselect		:IN		STD_LOGIC;
	avalon_read				:IN		STD_LOGIC;
	avalon_write			:IN		STD_LOGIC;
	avalon_writedata		:IN		STD_LOGIC_VECTOR(DW DOWNTO  0);	

	acknowledge				:IN		STD_LOGIC;
	irq						:IN		STD_LOGIC;
	read_data				:IN		STD_LOGIC_VECTOR(DW DOWNTO  0);	

	-- Bidirectionals

	-- Outputs
	avalon_irq				:BUFFER	STD_LOGIC;
	avalon_readdata		:BUFFER	STD_LOGIC_VECTOR(DW DOWNTO  0);	
	avalon_waitrequest	:BUFFER	STD_LOGIC;

	address					:BUFFER	STD_LOGIC_VECTOR(OW DOWNTO  0);	
	bus_enable				:BUFFER	STD_LOGIC;
	byte_enable				:BUFFER	STD_LOGIC_VECTOR(BW DOWNTO  0);	
	rw							:BUFFER	STD_LOGIC;
	write_data				:BUFFER	STD_LOGIC_VECTOR(DW DOWNTO  0)	

);

END nios_system_to_external_bus_bridge_0;

ARCHITECTURE Behaviour OF nios_system_to_external_bus_bridge_0 IS
-- *****************************************************************************
-- *                           Constant Declarations                           *
-- *****************************************************************************

-- *****************************************************************************
-- *                       Internal Signals Declarations                       *
-- *****************************************************************************
	
	-- Internal Wires
	
	-- Internal Registers
	SIGNAL	time_out_counter	:STD_LOGIC_VECTOR( 7 DOWNTO  0);	
	
	-- State Machine Registers
	
-- *****************************************************************************
-- *                          Component Declarations                           *
-- *****************************************************************************
BEGIN
-- *****************************************************************************
-- *                         Finite State Machine(s)                           *
-- *****************************************************************************


-- *****************************************************************************
-- *                             Sequential Logic                              *
-- *****************************************************************************

	PROCESS (clk)
	BEGIN
		IF clk'EVENT AND clk = '1' THEN
			IF (reset = '1') THEN
				avalon_readdata <= (OTHERS => '0');
			ELSIF ((acknowledge = '1') OR (AND_REDUCE(time_out_counter) = '1')) THEN
				avalon_readdata <= read_data;
			END IF;
		END IF;
	END PROCESS;


	PROCESS (clk)
	BEGIN
		IF clk'EVENT AND clk = '1' THEN
			IF (reset = '1') THEN
				address		<= (OTHERS => '0');
				bus_enable	<= '0';
				byte_enable	<= (OTHERS => '0');
				rw				<= '1';
				write_data	<= (OTHERS => '0');
			ELSE
				address		<= (avalon_address & (OTHERS => '0'));
		
				IF ((avalon_chipselect = '1') AND (OR_REDUCE(avalon_byteenable) = '1')) THEN
					bus_enable	<= avalon_waitrequest;
				ELSE
					bus_enable	<= '0';
		
			END IF;
				byte_enable	<= avalon_byteenable;
				rw				<= avalon_read OR NOT avalon_write;
				write_data	<= avalon_writedata;
			END IF;
		END IF;
	END PROCESS;


	PROCESS (clk)
	BEGIN
		IF clk'EVENT AND clk = '1' THEN
			IF (reset = '1') THEN
				time_out_counter <= B"00000000";
			ELSIF (avalon_waitrequest = '1') THEN
				time_out_counter <= time_out_counter + B"00000001";
			ELSE
				time_out_counter <= B"00000000";
			END IF;
		END IF;
	END PROCESS;


-- *****************************************************************************
-- *                            Combinational Logic                            *
-- *****************************************************************************

	avalon_irq 				<= irq;
	avalon_waitrequest 	<= 
			avalon_chipselect AND (OR_REDUCE(avalon_byteenable)) AND 
			 NOT acknowledge AND NOT (AND_REDUCE(time_out_counter));

-- *****************************************************************************
-- *                          Component Instantiations                         *
-- *****************************************************************************


END Behaviour;

